* Qucs 24.3.2  /home/denis/QucsWorkspace/voltage_devider_prj/main.sch
.INCLUDE "/tmp/.mount_Qucs-S6CkjU2/usr/share/qucs-s/xspice_cmlib/include/ngspice_mathfunc.inc"
V1 _net0 0 DC 100
R2 div2 _net1  1000 tc1=0.0 tc2=0.0 
R1 div1 _net2  455 tc1=0.0 tc2=0.0 
VPr1 _net0 _net2 DC 0
R6 0 _net3  5K tc1=0.0 tc2=0.0 
R5 _net4 0  2.5K tc1=0.0 tc2=0.0 
R7 0 _net5  2.5K tc1=0.0 tc2=0.0 
R4 0 _net6  5000 tc1=0.0 tc2=0.0 
VPr4 div3 _net6 DC 0
VPr2 div1 _net1 DC 0
VPr3 div2 _net7 DC 0
R3 div3 _net7  1680 tc1=0.0 tc2=0.0 
VPr5 div1 _net4 DC 0
VPr6 div2 _net3 DC 0
VPr7 div3 _net5 DC 0

.control

op
print i(VPr1) i(VPr2) i(VPr3) i(VPr4) i(VPr5) i(VPr6) i(VPr7) v(div1) v(div2) v(div3)   > spice4qucs.dc1.ngspice.dc.print
destroy all
reset

exit
.endc
.END
